module blockBottom(block, bottomY);

	input [0:8] block;
	output wire [1:0] bottomY;
	
	reg [0:8] tempBlock;
	reg [3:0] zeroNum;
	reg zeroStopFlag;
	reg [1:0] tempBottomY;
	integer i;
	
	always @(block) begin
		tempBlock = block; // Must be blocking assignment.
		zeroNum = 4'b0;
		zeroStopFlag = 1'b0;
		for (i = 0; i < 9; i = i + 1) begin
			if (tempBlock[8] == 1'b1) zeroStopFlag = 1'b1;
			else /*(tempBlock[8] == 1'b0)*/ begin
				zeroNum = zeroNum + 4'b1;
				//if (!zeroStopFlag) zeroNum = zeroNum + 4'b1;
				tempBlock = tempBlock >> 1'b1;
			end
		end
	end
	
	assign bottomY = zeroNum / 'd3;

endmodule
