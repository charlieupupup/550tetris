module background_always(
  input wire clk,
  input wire rst,
  input wire require_new_block, //1'b1 means the block is collided.
  input wire [4:0] blockX,
  input wire [4:0] blockY,

  input wire [15:0] block_rev,// 4*4 matrix

  output reg [399:0] field_display_out, //20*20 new background
  output wire [9:0] total_line_num
);

reg [9:0] total_line_num_inner;

wire [19:0] line; //representing whether each single line is full
wire is_any_line_full;

genvar gv_i;
generate for(gv_i = 0; gv_i < 20; gv_i = gv_i + 1)
    begin: line_check
        assign line[gv_i] = & field_display_out[(20 * gv_i + 19):(20 * gv_i)];
    end
endgenerate

assign is_any_line_full = | line[19:0]; //"is_any_line_full" is 1'd1 when at lease one line is full

initial begin
field_display_out <= 400'd0;
end

always @(posedge clk) begin
     if(is_any_line_full) begin
        if(line[0]) begin
            field_display_out[19:0]     <= 20'd0;
            field_display_out[39:20]    <= field_display_out[39:20]  ;
            field_display_out[59:40]    <= field_display_out[59:40]  ;
            field_display_out[79:60]    <= field_display_out[79:60]  ;
            field_display_out[99:80]    <= field_display_out[99:80]  ;
            field_display_out[119:100]  <= field_display_out[119:100];
            field_display_out[139:120]  <= field_display_out[139:120];
            field_display_out[159:140]  <= field_display_out[159:140];
            field_display_out[179:160]  <= field_display_out[179:160];
            field_display_out[199:180]  <= field_display_out[199:180];
            field_display_out[219:200]  <= field_display_out[219:200];
            field_display_out[239:220]  <= field_display_out[239:220];
            field_display_out[259:240]  <= field_display_out[259:240];
            field_display_out[279:260]  <= field_display_out[279:260];
            field_display_out[299:280]  <= field_display_out[299:280];
            field_display_out[319:300]  <= field_display_out[319:300];
            field_display_out[339:320]  <= field_display_out[339:320];
            field_display_out[359:340]  <= field_display_out[359:340];
            field_display_out[379:360]  <= field_display_out[379:360];
            field_display_out[399:380]  <= field_display_out[399:380];

            total_line_num_inner <= total_line_num_inner + 1; //full line recorder
        end

        if(line[1]) begin
            field_display_out[19:0]     <= 20'd0;
            field_display_out[39:20]    <= field_display_out[19:0]   ;
            field_display_out[59:40]    <= field_display_out[59:40]  ;
            field_display_out[79:60]    <= field_display_out[79:60]  ;
            field_display_out[99:80]    <= field_display_out[99:80]  ;
            field_display_out[119:100]  <= field_display_out[119:100];
            field_display_out[139:120]  <= field_display_out[139:120];
            field_display_out[159:140]  <= field_display_out[159:140];
            field_display_out[179:160]  <= field_display_out[179:160];
            field_display_out[199:180]  <= field_display_out[199:180];
            field_display_out[219:200]  <= field_display_out[219:200];
            field_display_out[239:220]  <= field_display_out[239:220];
            field_display_out[259:240]  <= field_display_out[259:240];
            field_display_out[279:260]  <= field_display_out[279:260];
            field_display_out[299:280]  <= field_display_out[299:280];
            field_display_out[319:300]  <= field_display_out[319:300];
            field_display_out[339:320]  <= field_display_out[339:320];
            field_display_out[359:340]  <= field_display_out[359:340];
            field_display_out[379:360]  <= field_display_out[379:360];
            field_display_out[399:380]  <= field_display_out[399:380];

            total_line_num_inner <= total_line_num_inner + 1; //full line recorder
        end

        if(line[2]) begin
            field_display_out[19:0]     <= 20'd0;
            field_display_out[39:20]    <= field_display_out[19:0]   ;
            field_display_out[59:40]    <= field_display_out[39:20]  ;
            field_display_out[79:60]    <= field_display_out[79:60]  ;
            field_display_out[99:80]    <= field_display_out[99:80]  ;
            field_display_out[119:100]  <= field_display_out[119:100];
            field_display_out[139:120]  <= field_display_out[139:120];
            field_display_out[159:140]  <= field_display_out[159:140];
            field_display_out[179:160]  <= field_display_out[179:160];
            field_display_out[199:180]  <= field_display_out[199:180];
            field_display_out[219:200]  <= field_display_out[219:200];
            field_display_out[239:220]  <= field_display_out[239:220];
            field_display_out[259:240]  <= field_display_out[259:240];
            field_display_out[279:260]  <= field_display_out[279:260];
            field_display_out[299:280]  <= field_display_out[299:280];
            field_display_out[319:300]  <= field_display_out[319:300];
            field_display_out[339:320]  <= field_display_out[339:320];
            field_display_out[359:340]  <= field_display_out[359:340];
            field_display_out[379:360]  <= field_display_out[379:360];
            field_display_out[399:380]  <= field_display_out[399:380];

            total_line_num_inner <= total_line_num_inner + 1; //full line recorder
        end

        if(line[3]) begin
            field_display_out[19:0]     <= 20'd0;
            field_display_out[39:20]    <= field_display_out[19:0]   ;
            field_display_out[59:40]    <= field_display_out[39:20]  ;
            field_display_out[79:60]    <= field_display_out[59:40]  ;
            field_display_out[99:80]    <= field_display_out[99:80]  ;
            field_display_out[119:100]  <= field_display_out[119:100];
            field_display_out[139:120]  <= field_display_out[139:120];
            field_display_out[159:140]  <= field_display_out[159:140];
            field_display_out[179:160]  <= field_display_out[179:160];
            field_display_out[199:180]  <= field_display_out[199:180];
            field_display_out[219:200]  <= field_display_out[219:200];
            field_display_out[239:220]  <= field_display_out[239:220];
            field_display_out[259:240]  <= field_display_out[259:240];
            field_display_out[279:260]  <= field_display_out[279:260];
            field_display_out[299:280]  <= field_display_out[299:280];
            field_display_out[319:300]  <= field_display_out[319:300];
            field_display_out[339:320]  <= field_display_out[339:320];
            field_display_out[359:340]  <= field_display_out[359:340];
            field_display_out[379:360]  <= field_display_out[379:360];
            field_display_out[399:380]  <= field_display_out[399:380];

            total_line_num_inner <= total_line_num_inner + 1; //full line recorder
        end

        if(line[4]) begin
            field_display_out[19:0]     <= 20'd0;
            field_display_out[39:20]    <= field_display_out[19:0]   ;
            field_display_out[59:40]    <= field_display_out[39:20]  ;
            field_display_out[79:60]    <= field_display_out[59:40]  ;
            field_display_out[99:80]    <= field_display_out[79:60]  ;
            field_display_out[119:100]  <= field_display_out[119:100];
            field_display_out[139:120]  <= field_display_out[139:120];
            field_display_out[159:140]  <= field_display_out[159:140];
            field_display_out[179:160]  <= field_display_out[179:160];
            field_display_out[199:180]  <= field_display_out[199:180];
            field_display_out[219:200]  <= field_display_out[219:200];
            field_display_out[239:220]  <= field_display_out[239:220];
            field_display_out[259:240]  <= field_display_out[259:240];
            field_display_out[279:260]  <= field_display_out[279:260];
            field_display_out[299:280]  <= field_display_out[299:280];
            field_display_out[319:300]  <= field_display_out[319:300];
            field_display_out[339:320]  <= field_display_out[339:320];
            field_display_out[359:340]  <= field_display_out[359:340];
            field_display_out[379:360]  <= field_display_out[379:360];
            field_display_out[399:380]  <= field_display_out[399:380];

            total_line_num_inner <= total_line_num_inner + 1; //full line recorder
        end

        if(line[5]) begin
            field_display_out[19:0]     <= 20'd0;
            field_display_out[39:20]    <= field_display_out[19:0]   ;
            field_display_out[59:40]    <= field_display_out[39:20]  ;
            field_display_out[79:60]    <= field_display_out[59:40]  ;
            field_display_out[99:80]    <= field_display_out[79:60]  ;
            field_display_out[119:100]  <= field_display_out[99:80]  ;
            field_display_out[139:120]  <= field_display_out[139:120];
            field_display_out[159:140]  <= field_display_out[159:140];
            field_display_out[179:160]  <= field_display_out[179:160];
            field_display_out[199:180]  <= field_display_out[199:180];
            field_display_out[219:200]  <= field_display_out[219:200];
            field_display_out[239:220]  <= field_display_out[239:220];
            field_display_out[259:240]  <= field_display_out[259:240];
            field_display_out[279:260]  <= field_display_out[279:260];
            field_display_out[299:280]  <= field_display_out[299:280];
            field_display_out[319:300]  <= field_display_out[319:300];
            field_display_out[339:320]  <= field_display_out[339:320];
            field_display_out[359:340]  <= field_display_out[359:340];
            field_display_out[379:360]  <= field_display_out[379:360];
            field_display_out[399:380]  <= field_display_out[399:380];

            total_line_num_inner <= total_line_num_inner + 1; //full line recorder
        end

        if(line[6]) begin
            field_display_out[19:0]     <= 20'd0;
            field_display_out[39:20]    <= field_display_out[19:0]   ;
            field_display_out[59:40]    <= field_display_out[39:20]  ;
            field_display_out[79:60]    <= field_display_out[59:40]  ;
            field_display_out[99:80]    <= field_display_out[79:60]  ;
            field_display_out[119:100]  <= field_display_out[99:80]  ;
            field_display_out[139:120]  <= field_display_out[119:100];
            field_display_out[159:140]  <= field_display_out[159:140];
            field_display_out[179:160]  <= field_display_out[179:160];
            field_display_out[199:180]  <= field_display_out[199:180];
            field_display_out[219:200]  <= field_display_out[219:200];
            field_display_out[239:220]  <= field_display_out[239:220];
            field_display_out[259:240]  <= field_display_out[259:240];
            field_display_out[279:260]  <= field_display_out[279:260];
            field_display_out[299:280]  <= field_display_out[299:280];
            field_display_out[319:300]  <= field_display_out[319:300];
            field_display_out[339:320]  <= field_display_out[339:320];
            field_display_out[359:340]  <= field_display_out[359:340];
            field_display_out[379:360]  <= field_display_out[379:360];
            field_display_out[399:380]  <= field_display_out[399:380];

            total_line_num_inner <= total_line_num_inner + 1; //full line recorder
        end

        if(line[7]) begin
            field_display_out[19:0]     <= 20'd0;
            field_display_out[39:20]    <= field_display_out[19:0]   ;
            field_display_out[59:40]    <= field_display_out[39:20]  ;
            field_display_out[79:60]    <= field_display_out[59:40]  ;
            field_display_out[99:80]    <= field_display_out[79:60]  ;
            field_display_out[119:100]  <= field_display_out[99:80]  ;
            field_display_out[139:120]  <= field_display_out[119:100];
            field_display_out[159:140]  <= field_display_out[139:120];
            field_display_out[179:160]  <= field_display_out[179:160];
            field_display_out[199:180]  <= field_display_out[199:180];
            field_display_out[219:200]  <= field_display_out[219:200];
            field_display_out[239:220]  <= field_display_out[239:220];
            field_display_out[259:240]  <= field_display_out[259:240];
            field_display_out[279:260]  <= field_display_out[279:260];
            field_display_out[299:280]  <= field_display_out[299:280];
            field_display_out[319:300]  <= field_display_out[319:300];
            field_display_out[339:320]  <= field_display_out[339:320];
            field_display_out[359:340]  <= field_display_out[359:340];
            field_display_out[379:360]  <= field_display_out[379:360];
            field_display_out[399:380]  <= field_display_out[399:380];

            total_line_num_inner <= total_line_num_inner + 1; //full line recorder
        end

        if(line[8]) begin
            field_display_out[19:0]     <= 20'd0;
            field_display_out[39:20]    <= field_display_out[19:0]   ;
            field_display_out[59:40]    <= field_display_out[39:20]  ;
            field_display_out[79:60]    <= field_display_out[59:40]  ;
            field_display_out[99:80]    <= field_display_out[79:60]  ;
            field_display_out[119:100]  <= field_display_out[99:80]  ;
            field_display_out[139:120]  <= field_display_out[119:100];
            field_display_out[159:140]  <= field_display_out[139:120];
            field_display_out[179:160]  <= field_display_out[159:140];
            field_display_out[199:180]  <= field_display_out[199:180];
            field_display_out[219:200]  <= field_display_out[219:200];
            field_display_out[239:220]  <= field_display_out[239:220];
            field_display_out[259:240]  <= field_display_out[259:240];
            field_display_out[279:260]  <= field_display_out[279:260];
            field_display_out[299:280]  <= field_display_out[299:280];
            field_display_out[319:300]  <= field_display_out[319:300];
            field_display_out[339:320]  <= field_display_out[339:320];
            field_display_out[359:340]  <= field_display_out[359:340];
            field_display_out[379:360]  <= field_display_out[379:360];
            field_display_out[399:380]  <= field_display_out[399:380];

            total_line_num_inner <= total_line_num_inner + 1; //full line recorder
        end

        if(line[9]) begin
            field_display_out[19:0]     <= 20'd0;
            field_display_out[39:20]    <= field_display_out[19:0]   ;
            field_display_out[59:40]    <= field_display_out[39:20]  ;
            field_display_out[79:60]    <= field_display_out[59:40]  ;
            field_display_out[99:80]    <= field_display_out[79:60]  ;
            field_display_out[119:100]  <= field_display_out[99:80]  ;
            field_display_out[139:120]  <= field_display_out[119:100];
            field_display_out[159:140]  <= field_display_out[139:120];
            field_display_out[179:160]  <= field_display_out[159:140];
            field_display_out[199:180]  <= field_display_out[179:160];
            field_display_out[219:200]  <= field_display_out[219:200];
            field_display_out[239:220]  <= field_display_out[239:220];
            field_display_out[259:240]  <= field_display_out[259:240];
            field_display_out[279:260]  <= field_display_out[279:260];
            field_display_out[299:280]  <= field_display_out[299:280];
            field_display_out[319:300]  <= field_display_out[319:300];
            field_display_out[339:320]  <= field_display_out[339:320];
            field_display_out[359:340]  <= field_display_out[359:340];
            field_display_out[379:360]  <= field_display_out[379:360];
            field_display_out[399:380]  <= field_display_out[399:380];

            total_line_num_inner <= total_line_num_inner + 1; //full line recorder
        end

        if(line[10]) begin
            field_display_out[19:0]     <= 20'd0;
            field_display_out[39:20]    <= field_display_out[19:0]   ;
            field_display_out[59:40]    <= field_display_out[39:20]  ;
            field_display_out[79:60]    <= field_display_out[59:40]  ;
            field_display_out[99:80]    <= field_display_out[79:60]  ;
            field_display_out[119:100]  <= field_display_out[99:80]  ;
            field_display_out[139:120]  <= field_display_out[119:100];
            field_display_out[159:140]  <= field_display_out[139:120];
            field_display_out[179:160]  <= field_display_out[159:140];
            field_display_out[199:180]  <= field_display_out[179:160];
            field_display_out[219:200]  <= field_display_out[199:180];
            field_display_out[239:220]  <= field_display_out[239:220];
            field_display_out[259:240]  <= field_display_out[259:240];
            field_display_out[279:260]  <= field_display_out[279:260];
            field_display_out[299:280]  <= field_display_out[299:280];
            field_display_out[319:300]  <= field_display_out[319:300];
            field_display_out[339:320]  <= field_display_out[339:320];
            field_display_out[359:340]  <= field_display_out[359:340];
            field_display_out[379:360]  <= field_display_out[379:360];
            field_display_out[399:380]  <= field_display_out[399:380];

            total_line_num_inner <= total_line_num_inner + 1; //full line recorder
        end

        if(line[11]) begin
            field_display_out[19:0]     <= 20'd0;
            field_display_out[39:20]    <= field_display_out[19:0]   ;
            field_display_out[59:40]    <= field_display_out[39:20]  ;
            field_display_out[79:60]    <= field_display_out[59:40]  ;
            field_display_out[99:80]    <= field_display_out[79:60]  ;
            field_display_out[119:100]  <= field_display_out[99:80]  ;
            field_display_out[139:120]  <= field_display_out[119:100];
            field_display_out[159:140]  <= field_display_out[139:120];
            field_display_out[179:160]  <= field_display_out[159:140];
            field_display_out[199:180]  <= field_display_out[179:160];
            field_display_out[219:200]  <= field_display_out[199:180];
            field_display_out[239:220]  <= field_display_out[219:200];
            field_display_out[259:240]  <= field_display_out[259:240];
            field_display_out[279:260]  <= field_display_out[279:260];
            field_display_out[299:280]  <= field_display_out[299:280];
            field_display_out[319:300]  <= field_display_out[319:300];
            field_display_out[339:320]  <= field_display_out[339:320];
            field_display_out[359:340]  <= field_display_out[359:340];
            field_display_out[379:360]  <= field_display_out[379:360];
            field_display_out[399:380]  <= field_display_out[399:380];

            total_line_num_inner <= total_line_num_inner + 1; //full line recorder
        end

        if(line[12]) begin
            field_display_out[19:0]     <= 20'd0;
            field_display_out[39:20]    <= field_display_out[19:0]   ;
            field_display_out[59:40]    <= field_display_out[39:20]  ;
            field_display_out[79:60]    <= field_display_out[59:40]  ;
            field_display_out[99:80]    <= field_display_out[79:60]  ;
            field_display_out[119:100]  <= field_display_out[99:80]  ;
            field_display_out[139:120]  <= field_display_out[119:100];
            field_display_out[159:140]  <= field_display_out[139:120];
            field_display_out[179:160]  <= field_display_out[159:140];
            field_display_out[199:180]  <= field_display_out[179:160];
            field_display_out[219:200]  <= field_display_out[199:180];
            field_display_out[239:220]  <= field_display_out[219:200];
            field_display_out[259:240]  <= field_display_out[239:220];
            field_display_out[279:260]  <= field_display_out[279:260];
            field_display_out[299:280]  <= field_display_out[299:280];
            field_display_out[319:300]  <= field_display_out[319:300];
            field_display_out[339:320]  <= field_display_out[339:320];
            field_display_out[359:340]  <= field_display_out[359:340];
            field_display_out[379:360]  <= field_display_out[379:360];
            field_display_out[399:380]  <= field_display_out[399:380];

            total_line_num_inner <= total_line_num_inner + 1; //full line recorder
        end

        if(line[13]) begin
            field_display_out[19:0]     <= 20'd0;
            field_display_out[39:20]    <= field_display_out[19:0]   ;
            field_display_out[59:40]    <= field_display_out[39:20]  ;
            field_display_out[79:60]    <= field_display_out[59:40]  ;
            field_display_out[99:80]    <= field_display_out[79:60]  ;
            field_display_out[119:100]  <= field_display_out[99:80]  ;
            field_display_out[139:120]  <= field_display_out[119:100];
            field_display_out[159:140]  <= field_display_out[139:120];
            field_display_out[179:160]  <= field_display_out[159:140];
            field_display_out[199:180]  <= field_display_out[179:160];
            field_display_out[219:200]  <= field_display_out[199:180];
            field_display_out[239:220]  <= field_display_out[219:200];
            field_display_out[259:240]  <= field_display_out[239:220];
            field_display_out[279:260]  <= field_display_out[259:240];
            field_display_out[299:280]  <= field_display_out[299:280];
            field_display_out[319:300]  <= field_display_out[319:300];
            field_display_out[339:320]  <= field_display_out[339:320];
            field_display_out[359:340]  <= field_display_out[359:340];
            field_display_out[379:360]  <= field_display_out[379:360];
            field_display_out[399:380]  <= field_display_out[399:380];

            total_line_num_inner <= total_line_num_inner + 1; //full line recorder
        end

        if(line[14]) begin
            field_display_out[19:0]     <= 20'd0;
            field_display_out[39:20]    <= field_display_out[19:0]   ;
            field_display_out[59:40]    <= field_display_out[39:20]  ;
            field_display_out[79:60]    <= field_display_out[59:40]  ;
            field_display_out[99:80]    <= field_display_out[79:60]  ;
            field_display_out[119:100]  <= field_display_out[99:80]  ;
            field_display_out[139:120]  <= field_display_out[119:100];
            field_display_out[159:140]  <= field_display_out[139:120];
            field_display_out[179:160]  <= field_display_out[159:140];
            field_display_out[199:180]  <= field_display_out[179:160];
            field_display_out[219:200]  <= field_display_out[199:180];
            field_display_out[239:220]  <= field_display_out[219:200];
            field_display_out[259:240]  <= field_display_out[239:220];
            field_display_out[279:260]  <= field_display_out[259:240];
            field_display_out[299:280]  <= field_display_out[279:260];
            field_display_out[319:300]  <= field_display_out[319:300];
            field_display_out[339:320]  <= field_display_out[339:320];
            field_display_out[359:340]  <= field_display_out[359:340];
            field_display_out[379:360]  <= field_display_out[379:360];
            field_display_out[399:380]  <= field_display_out[399:380];

            total_line_num_inner <= total_line_num_inner + 1; //full line recorder
        end

        if(line[15]) begin
            field_display_out[19:0]     <= 20'd0;
            field_display_out[39:20]    <= field_display_out[19:0]   ;
            field_display_out[59:40]    <= field_display_out[39:20]  ;
            field_display_out[79:60]    <= field_display_out[59:40]  ;
            field_display_out[99:80]    <= field_display_out[79:60]  ;
            field_display_out[119:100]  <= field_display_out[99:80]  ;
            field_display_out[139:120]  <= field_display_out[119:100];
            field_display_out[159:140]  <= field_display_out[139:120];
            field_display_out[179:160]  <= field_display_out[159:140];
            field_display_out[199:180]  <= field_display_out[179:160];
            field_display_out[219:200]  <= field_display_out[199:180];
            field_display_out[239:220]  <= field_display_out[219:200];
            field_display_out[259:240]  <= field_display_out[239:220];
            field_display_out[279:260]  <= field_display_out[259:240];
            field_display_out[299:280]  <= field_display_out[279:260];
            field_display_out[319:300]  <= field_display_out[299:280];
            field_display_out[339:320]  <= field_display_out[339:320];
            field_display_out[359:340]  <= field_display_out[359:340];
            field_display_out[379:360]  <= field_display_out[379:360];
            field_display_out[399:380]  <= field_display_out[399:380];

            total_line_num_inner <= total_line_num_inner + 1; //full line recorder
        end

        if(line[16]) begin
            field_display_out[19:0]     <= 20'd0;
            field_display_out[39:20]    <= field_display_out[19:0]   ;
            field_display_out[59:40]    <= field_display_out[39:20]  ;
            field_display_out[79:60]    <= field_display_out[59:40]  ;
            field_display_out[99:80]    <= field_display_out[79:60]  ;
            field_display_out[119:100]  <= field_display_out[99:80]  ;
            field_display_out[139:120]  <= field_display_out[119:100];
            field_display_out[159:140]  <= field_display_out[139:120];
            field_display_out[179:160]  <= field_display_out[159:140];
            field_display_out[199:180]  <= field_display_out[179:160];
            field_display_out[219:200]  <= field_display_out[199:180];
            field_display_out[239:220]  <= field_display_out[219:200];
            field_display_out[259:240]  <= field_display_out[239:220];
            field_display_out[279:260]  <= field_display_out[259:240];
            field_display_out[299:280]  <= field_display_out[279:260];
            field_display_out[319:300]  <= field_display_out[299:280];
            field_display_out[339:320]  <= field_display_out[319:300];
            field_display_out[359:340]  <= field_display_out[359:340];
            field_display_out[379:360]  <= field_display_out[379:360];
            field_display_out[399:380]  <= field_display_out[399:380];

            total_line_num_inner <= total_line_num_inner + 1; //full line recorder
        end

        if(line[17]) begin
            field_display_out[19:0]     <= 20'd0;
            field_display_out[39:20]    <= field_display_out[19:0]   ;
            field_display_out[59:40]    <= field_display_out[39:20]  ;
            field_display_out[79:60]    <= field_display_out[59:40]  ;
            field_display_out[99:80]    <= field_display_out[79:60]  ;
            field_display_out[119:100]  <= field_display_out[99:80]  ;
            field_display_out[139:120]  <= field_display_out[119:100];
            field_display_out[159:140]  <= field_display_out[139:120];
            field_display_out[179:160]  <= field_display_out[159:140];
            field_display_out[199:180]  <= field_display_out[179:160];
            field_display_out[219:200]  <= field_display_out[199:180];
            field_display_out[239:220]  <= field_display_out[219:200];
            field_display_out[259:240]  <= field_display_out[239:220];
            field_display_out[279:260]  <= field_display_out[259:240];
            field_display_out[299:280]  <= field_display_out[279:260];
            field_display_out[319:300]  <= field_display_out[299:280];
            field_display_out[339:320]  <= field_display_out[319:300];
            field_display_out[359:340]  <= field_display_out[339:320];
            field_display_out[379:360]  <= field_display_out[379:360];
            field_display_out[399:380]  <= field_display_out[399:380];

            total_line_num_inner <= total_line_num_inner + 1; //full line recorder
        end

        if(line[18]) begin
            field_display_out[19:0]     <= 20'd0;
            field_display_out[39:20]    <= field_display_out[19:0]   ;
            field_display_out[59:40]    <= field_display_out[39:20]  ;
            field_display_out[79:60]    <= field_display_out[59:40]  ;
            field_display_out[99:80]    <= field_display_out[79:60]  ;
            field_display_out[119:100]  <= field_display_out[99:80]  ;
            field_display_out[139:120]  <= field_display_out[119:100];
            field_display_out[159:140]  <= field_display_out[139:120];
            field_display_out[179:160]  <= field_display_out[159:140];
            field_display_out[199:180]  <= field_display_out[179:160];
            field_display_out[219:200]  <= field_display_out[199:180];
            field_display_out[239:220]  <= field_display_out[219:200];
            field_display_out[259:240]  <= field_display_out[239:220];
            field_display_out[279:260]  <= field_display_out[259:240];
            field_display_out[299:280]  <= field_display_out[279:260];
            field_display_out[319:300]  <= field_display_out[299:280];
            field_display_out[339:320]  <= field_display_out[319:300];
            field_display_out[359:340]  <= field_display_out[339:320];
            field_display_out[379:360]  <= field_display_out[359:340];
            field_display_out[399:380]  <= field_display_out[399:380];

            total_line_num_inner <= total_line_num_inner + 1; //full line recorder
        end

        if(line[19]) begin
            field_display_out[19:0]     <= 20'd0;
            field_display_out[39:20]    <= field_display_out[19:0]   ;
            field_display_out[59:40]    <= field_display_out[39:20]  ;
            field_display_out[79:60]    <= field_display_out[59:40]  ;
            field_display_out[99:80]    <= field_display_out[79:60]  ;
            field_display_out[119:100]  <= field_display_out[99:80]  ;
            field_display_out[139:120]  <= field_display_out[119:100];
            field_display_out[159:140]  <= field_display_out[139:120];
            field_display_out[179:160]  <= field_display_out[159:140];
            field_display_out[199:180]  <= field_display_out[179:160];
            field_display_out[219:200]  <= field_display_out[199:180];
            field_display_out[239:220]  <= field_display_out[219:200];
            field_display_out[259:240]  <= field_display_out[239:220];
            field_display_out[279:260]  <= field_display_out[259:240];
            field_display_out[299:280]  <= field_display_out[279:260];
            field_display_out[319:300]  <= field_display_out[299:280];
            field_display_out[339:320]  <= field_display_out[319:300];
            field_display_out[359:340]  <= field_display_out[339:320];
            field_display_out[379:360]  <= field_display_out[359:340];
            field_display_out[399:380]  <= field_display_out[379:360];

            total_line_num_inner <= total_line_num_inner + 1; //full line recorder
        end
    end

    else if( require_new_block ) begin
        field_display_out[blockY * 20 + blockX + 5'd0] <= block_rev[0] || field_display_out[blockY * 20 + blockX + 5'd0];
        field_display_out[blockY * 20 + blockX + 5'd1] <= block_rev[1] || field_display_out[blockY * 20 + blockX + 5'd1];
        field_display_out[blockY * 20 + blockX + 5'd2] <= block_rev[2] || field_display_out[blockY * 20 + blockX + 5'd2];
        field_display_out[blockY * 20 + blockX + 5'd3] <= block_rev[3] || field_display_out[blockY * 20 + blockX + 5'd3];        
        field_display_out[blockY * 20 + blockX + 5'd20] <= block_rev[4] || field_display_out[blockY * 20 + blockX + 5'd20];
        field_display_out[blockY * 20 + blockX + 5'd21] <= block_rev[5] || field_display_out[blockY * 20 + blockX + 5'd21];
        field_display_out[blockY * 20 + blockX + 5'd22] <= block_rev[6] || field_display_out[blockY * 20 + blockX + 5'd22];
        field_display_out[blockY * 20 + blockX + 5'd23] <= block_rev[7] || field_display_out[blockY * 20 + blockX + 5'd23];    
        field_display_out[blockY * 20 + blockX + 5'd40] <= block_rev[8] || field_display_out[blockY * 20 + blockX + 5'd40];
        field_display_out[blockY * 20 + blockX + 5'd41] <= block_rev[9] || field_display_out[blockY * 20 + blockX + 5'd41];
        field_display_out[blockY * 20 + blockX + 5'd42] <= block_rev[10] || field_display_out[blockY * 20 + blockX + 5'd42];
        field_display_out[blockY * 20 + blockX + 5'd43] <= block_rev[11] || field_display_out[blockY * 20 + blockX + 5'd43];        
        field_display_out[blockY * 20 + blockX + 5'd60] <= block_rev[12] || field_display_out[blockY * 20 + blockX + 5'd60];
        field_display_out[blockY * 20 + blockX + 5'd61] <= block_rev[13] || field_display_out[blockY * 20 + blockX + 5'd61];
        field_display_out[blockY * 20 + blockX + 5'd62] <= block_rev[14] || field_display_out[blockY * 20 + blockX + 5'd62];
        field_display_out[blockY * 20 + blockX + 5'd63] <= block_rev[15] || field_display_out[blockY * 20 + blockX + 5'd63];
        total_line_num_inner <= total_line_num_inner ;
      end
		end

  assign total_line_num = total_line_num_inner;
    


endmodule
